
/*****************************************************************************************************
 * Copyright (c) 2024 SiPlusPlus Semiconductor
 *
 * FileContributor: Dinesh Annayya <dinesha@opencores.org>                       
 * FileContributor: Dinesh Annayya <dinesh@siplusplus.com>                       
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *      http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 ***************************************************************************************************/
`ifndef CACHE_INCLUDE_DEFS
`define CACHE_INCLUDE_DEFS

`define TAG_XLEN        20

// Tag Memory List
typedef struct packed {
    logic                             valid;
    logic                             dirty;
    logic [`TAG_XLEN-1:0]             tag;
} type_dcache_tag_mem_s;

// Tag Memory List
typedef struct packed {
    logic                             valid;
    logic [`TAG_XLEN-1:0]             tag;
} type_icache_tag_mem_s;

`endif
